--==============================================================================
--== Logisim goes FPGA automatic generated VHDL code                          ==
--==                                                                          ==
--==                                                                          ==
--== Project   : exampleLog                                                   ==
--== Component : main                                                         ==
--==                                                                          ==
--==============================================================================


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY main IS
   PORT ( asd                       : IN  std_logic;
          bsd                       : IN  std_logic;
          ccs                       : OUT std_logic);
END main;

