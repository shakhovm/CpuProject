--==============================================================================
--== Logisim goes FPGA automatic generated VHDL code                          ==
--==                                                                          ==
--==                                                                          ==
--== Project   : exampleLog                                                   ==
--== Component : LogisimToplevelShell                                         ==
--==                                                                          ==
--==============================================================================


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY LogisimToplevelShell IS
   PORT ( FPGA_INPUT_PIN_0          : IN  std_logic;
          FPGA_INPUT_PIN_1          : IN  std_logic;
          FPGA_OUTPUT_PIN_0         : OUT std_logic);
END LogisimToplevelShell;

